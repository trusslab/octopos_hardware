`include "./Octopos_MailBox_Main_logic.v"
`include "./Octopos_MailBox_Ctrl_Interface_Manager.v"
`include "./Octopos_MailBox_ctrl_AXI.v"
`include "./Octopos_MailBox_1Writer_3Reader_v1_0.v"

module top
(
	// MailBox Main Signals
	input wire S_CLK,
	input wire S_ARESETN,
	// Ctrl0 AXI port
	input wire  s_ctrl0_axi_aclk,
	input wire  s_ctrl0_axi_aresetn,
	input wire [3 : 0] s_ctrl0_axi_awaddr,
	input wire [2 : 0] s_ctrl0_axi_awprot,
	input wire  s_ctrl0_axi_awvalid,
	output wire  s_ctrl0_axi_awready,
	input wire [31 : 0] s_ctrl0_axi_wdata,
	input wire [3 : 0] s_ctrl0_axi_wstrb,
	input wire  s_ctrl0_axi_wvalid,
	output wire  s_ctrl0_axi_wready,
	output wire [1 : 0] s_ctrl0_axi_bresp,
	output wire  s_ctrl0_axi_bvalid,
	input wire  s_ctrl0_axi_bready,
	input wire [3 : 0] s_ctrl0_axi_araddr,
	input wire [2 : 0] s_ctrl0_axi_arprot,
	input wire  s_ctrl0_axi_arvalid,
	output wire  s_ctrl0_axi_arready,
	output wire [31 : 0] s_ctrl0_axi_rdata,
	output wire [1 : 0] s_ctrl0_axi_rresp,
	output wire  s_ctrl0_axi_rvalid,
	input wire  s_ctrl0_axi_rready,
	// Ctrl1 AXI port
	input wire  s_ctrl1_axi_aclk,
	input wire  s_ctrl1_axi_aresetn,
	input wire [3 : 0] s_ctrl1_axi_awaddr,
	input wire [2 : 0] s_ctrl1_axi_awprot,
	input wire  s_ctrl1_axi_awvalid,
	output wire  s_ctrl1_axi_awready,
	input wire [31 : 0] s_ctrl1_axi_wdata,
	input wire [3 : 0] s_ctrl1_axi_wstrb,
	input wire  s_ctrl1_axi_wvalid,
	output wire  s_ctrl1_axi_wready,
	output wire [1 : 0] s_ctrl1_axi_bresp,
	output wire  s_ctrl1_axi_bvalid,
	input wire  s_ctrl1_axi_bready,
	input wire [3 : 0] s_ctrl1_axi_araddr,
	input wire [2 : 0] s_ctrl1_axi_arprot,
	input wire  s_ctrl1_axi_arvalid,
	output wire  s_ctrl1_axi_arready,
	output wire [31 : 0] s_ctrl1_axi_rdata,
	output wire [1 : 0] s_ctrl1_axi_rresp,
	output wire  s_ctrl1_axi_rvalid,
	input wire  s_ctrl1_axi_rready,
	// Ctrl2 AXI port
	input wire  s_ctrl2_axi_aclk,
	input wire  s_ctrl2_axi_aresetn,
	input wire [3 : 0] s_ctrl2_axi_awaddr,
	input wire [2 : 0] s_ctrl2_axi_awprot,
	input wire  s_ctrl2_axi_awvalid,
	output wire  s_ctrl2_axi_awready,
	input wire [31 : 0] s_ctrl2_axi_wdata,
	input wire [3 : 0] s_ctrl2_axi_wstrb,
	input wire  s_ctrl2_axi_wvalid,
	output wire  s_ctrl2_axi_wready,
	output wire [1 : 0] s_ctrl2_axi_bresp,
	output wire  s_ctrl2_axi_bvalid,
	input wire  s_ctrl2_axi_bready,
	input wire [3 : 0] s_ctrl2_axi_araddr,
	input wire [2 : 0] s_ctrl2_axi_arprot,
	input wire  s_ctrl2_axi_arvalid,
	output wire  s_ctrl2_axi_arready,
	output wire [31 : 0] s_ctrl2_axi_rdata,
	output wire [1 : 0] s_ctrl2_axi_rresp,
	output wire  s_ctrl2_axi_rvalid,
	input wire  s_ctrl2_axi_rready,
	// Ctrl_fixed AXI port
	input wire  s_ctrl_fixed_axi_aclk,
	input wire  s_ctrl_fixed_axi_aresetn,
	input wire [3 : 0] s_ctrl_fixed_axi_awaddr,
	input wire [2 : 0] s_ctrl_fixed_axi_awprot,
	input wire  s_ctrl_fixed_axi_awvalid,
	output wire  s_ctrl_fixed_axi_awready,
	input wire [31 : 0] s_ctrl_fixed_axi_wdata,
	input wire [3 : 0] s_ctrl_fixed_axi_wstrb,
	input wire  s_ctrl_fixed_axi_wvalid,
	output wire  s_ctrl_fixed_axi_wready,
	output wire [1 : 0] s_ctrl_fixed_axi_bresp,
	output wire  s_ctrl_fixed_axi_bvalid,
	input wire  s_ctrl_fixed_axi_bready,
	input wire [3 : 0] s_ctrl_fixed_axi_araddr,
	input wire [2 : 0] s_ctrl_fixed_axi_arprot,
	input wire  s_ctrl_fixed_axi_arvalid,
	output wire  s_ctrl_fixed_axi_arready,
	output wire [31 : 0] s_ctrl_fixed_axi_rdata,
	output wire [1 : 0] s_ctrl_fixed_axi_rresp,
	output wire  s_ctrl_fixed_axi_rvalid,
	input wire  s_ctrl_fixed_axi_rready,
	// data0 AXI port
	input wire S0_data0_AXI_ACLK,
	input wire S0_data0_AXI_ARESETN,
	input wire [31 : 0] S0_data0_AXI_AWADDR,
	input wire S0_data0_AXI_AWVALID,
	output wire S0_data0_AXI_AWREADY,
	input wire [31 : 0] S0_data0_AXI_WDATA,
	input wire [3 : 0] S0_data0_AXI_WSTRB,
	input wire S0_data0_AXI_WVALID,
	output wire S0_data0_AXI_WREADY,
	output wire [1 : 0] S0_data0_AXI_BRESP,
	output wire S0_data0_AXI_BVALID,
	input wire S0_data0_AXI_BREADY,
	input wire [31 : 0] S0_data0_AXI_ARADDR,
	input wire S0_data0_AXI_ARVALID,
	output wire S0_data0_AXI_ARREADY,
	output wire [31 : 0] S0_data0_AXI_RDATA,
	output wire [1 : 0] S0_data0_AXI_RRESP,
	output wire S0_data0_AXI_RVALID,
	input wire S0_data0_AXI_RREADY,
	// data1 AXI port
	input wire S0_data1_AXI_ACLK,
	input wire S0_data1_AXI_ARESETN,
	input wire [31 : 0] S0_data1_AXI_AWADDR,
	input wire S0_data1_AXI_AWVALID,
	output wire S0_data1_AXI_AWREADY,
	input wire [31 : 0] S0_data1_AXI_WDATA,
	input wire [3 : 0] S0_data1_AXI_WSTRB,
	input wire S0_data1_AXI_WVALID,
	output wire S0_data1_AXI_WREADY,
	output wire [1 : 0] S0_data1_AXI_BRESP,
	output wire S0_data1_AXI_BVALID,
	input wire S0_data1_AXI_BREADY,
	input wire [31 : 0] S0_data1_AXI_ARADDR,
	input wire S0_data1_AXI_ARVALID,
	output wire S0_data1_AXI_ARREADY,
	output wire [31 : 0] S0_data1_AXI_RDATA,
	output wire [1 : 0] S0_data1_AXI_RRESP,
	output wire S0_data1_AXI_RVALID,
	input wire S0_data1_AXI_RREADY,
	// data2 AXI port
	input wire S0_data2_AXI_ACLK,
	input wire S0_data2_AXI_ARESETN,
	input wire [31 : 0] S0_data2_AXI_AWADDR,
	input wire S0_data2_AXI_AWVALID,
	output wire S0_data2_AXI_AWREADY,
	input wire [31 : 0] S0_data2_AXI_WDATA,
	input wire [3 : 0] S0_data2_AXI_WSTRB,
	input wire S0_data2_AXI_WVALID,
	output wire S0_data2_AXI_WREADY,
	output wire [1 : 0] S0_data2_AXI_BRESP,
	output wire S0_data2_AXI_BVALID,
	input wire S0_data2_AXI_BREADY,
	input wire [31 : 0] S0_data2_AXI_ARADDR,
	input wire S0_data2_AXI_ARVALID,
	output wire S0_data2_AXI_ARREADY,
	output wire [31 : 0] S0_data2_AXI_RDATA,
	output wire [1 : 0] S0_data2_AXI_RRESP,
	output wire S0_data2_AXI_RVALID,
	input wire S0_data2_AXI_RREADY,
	// data_fixed AXI port
	input wire S1_data_fixed_AXI_ACLK,
	input wire S1_data_fixed_AXI_ARESETN,
	input wire [31 : 0] S1_data_fixed_AXI_AWADDR,
	input wire S1_data_fixed_AXI_AWVALID,
	output wire S1_data_fixed_AXI_AWREADY,
	input wire [31 : 0] S1_data_fixed_AXI_WDATA,
	input wire [3 : 0] S1_data_fixed_AXI_WSTRB,
	input wire S1_data_fixed_AXI_WVALID,
	output wire S1_data_fixed_AXI_WREADY,
	output wire [1 : 0] S1_data_fixed_AXI_BRESP,
	output wire S1_data_fixed_AXI_BVALID,
	input wire S1_data_fixed_AXI_BREADY,
	input wire [31 : 0] S1_data_fixed_AXI_ARADDR,
	input wire S1_data_fixed_AXI_ARVALID,
	output wire S1_data_fixed_AXI_ARREADY,
	output wire [31 : 0] S1_data_fixed_AXI_RDATA,
	output wire [1 : 0] S1_data_fixed_AXI_RRESP,
	output wire S1_data_fixed_AXI_RVALID,
	input wire S1_data_fixed_AXI_RREADY,
	// Interrupt lines
	output wire Interrupt_0,
	output wire Interrupt_ctrl0,
	output wire Interrupt_1,
	output wire Interrupt_ctrl1,
	output wire Interrupt_2,
	output wire Interrupt_ctrl2,
	output wire Interrupt_fixed,
	output wire Interrupt_ctrl_fixed,
	output wire busy0,
	output wire busy1,
	output wire busy2,
	output wire busy3,
	output wire busy4,
	output wire busy5,
	output wire busy6,
	output wire busy7,
	//tmp output for verification
	output wire [31:0] state_reg_out,
	output wire [31:0] S0_data_AXI_WDATA,
	output wire [31:0] S0_data_AXI_RDATA

);//Ports def end


Octopos_MailBox_1Writer_3Reader_v1_0 uut (
	// MailBox Main Signals
	S_CLK,
	S_ARESETN,
	// Ctrl0 AXI port
	s_ctrl0_axi_aclk,
	s_ctrl0_axi_aresetn,
	s_ctrl0_axi_awaddr,
	s_ctrl0_axi_awprot,
	s_ctrl0_axi_awvalid,
	s_ctrl0_axi_awready,
	s_ctrl0_axi_wdata,
	s_ctrl0_axi_wstrb,
	s_ctrl0_axi_wvalid,
	s_ctrl0_axi_wready,
	s_ctrl0_axi_bresp,
	s_ctrl0_axi_bvalid,
	s_ctrl0_axi_bready,
	s_ctrl0_axi_araddr,
	s_ctrl0_axi_arprot,
	s_ctrl0_axi_arvalid,
	s_ctrl0_axi_arready,
	s_ctrl0_axi_rdata,
	s_ctrl0_axi_rresp,
	s_ctrl0_axi_rvalid,
	s_ctrl0_axi_rready,
	// Ctrl1 AXI port
	s_ctrl1_axi_aclk,
	s_ctrl1_axi_aresetn,
	s_ctrl1_axi_awaddr,
	s_ctrl1_axi_awprot,
	s_ctrl1_axi_awvalid,
	s_ctrl1_axi_awready,
	s_ctrl1_axi_wdata,
	s_ctrl1_axi_wstrb,
	s_ctrl1_axi_wvalid,
	s_ctrl1_axi_wready,
	s_ctrl1_axi_bresp,
	s_ctrl1_axi_bvalid,
	s_ctrl1_axi_bready,
	s_ctrl1_axi_araddr,
	s_ctrl1_axi_arprot,
	s_ctrl1_axi_arvalid,
	s_ctrl1_axi_arready,
	s_ctrl1_axi_rdata,
	s_ctrl1_axi_rresp,
	s_ctrl1_axi_rvalid,
	s_ctrl1_axi_rready,
	// Ctrl2 AXI port
	s_ctrl2_axi_aclk,
	s_ctrl2_axi_aresetn,
	s_ctrl2_axi_awaddr,
	s_ctrl2_axi_awprot,
	s_ctrl2_axi_awvalid,
	s_ctrl2_axi_awready,
	s_ctrl2_axi_wdata,
	s_ctrl2_axi_wstrb,
	s_ctrl2_axi_wvalid,
	s_ctrl2_axi_wready,
	s_ctrl2_axi_bresp,
	s_ctrl2_axi_bvalid,
	s_ctrl2_axi_bready,
	s_ctrl2_axi_araddr,
	s_ctrl2_axi_arprot,
	s_ctrl2_axi_arvalid,
	s_ctrl2_axi_arready,
	s_ctrl2_axi_rdata,
	s_ctrl2_axi_rresp,
	s_ctrl2_axi_rvalid,
	s_ctrl2_axi_rready,
	// Ctrl_fixed AXI port
	s_ctrl_fixed_axi_aclk,
	s_ctrl_fixed_axi_aresetn,
	s_ctrl_fixed_axi_awaddr,
	s_ctrl_fixed_axi_awprot,
	s_ctrl_fixed_axi_awvalid,
	s_ctrl_fixed_axi_awready,
	s_ctrl_fixed_axi_wdata,
	s_ctrl_fixed_axi_wstrb,
	s_ctrl_fixed_axi_wvalid,
	s_ctrl_fixed_axi_wready,
	s_ctrl_fixed_axi_bresp,
	s_ctrl_fixed_axi_bvalid,
	s_ctrl_fixed_axi_bready,
	s_ctrl_fixed_axi_araddr,
	s_ctrl_fixed_axi_arprot,
	s_ctrl_fixed_axi_arvalid,
	s_ctrl_fixed_axi_arready,
	s_ctrl_fixed_axi_rdata,
	s_ctrl_fixed_axi_rresp,
	s_ctrl_fixed_axi_rvalid,
	s_ctrl_fixed_axi_rready,
	// data0 AXI port
	S0_data0_AXI_ACLK,
	S0_data0_AXI_ARESETN,
	S0_data0_AXI_AWADDR,
	S0_data0_AXI_AWVALID,
	S0_data0_AXI_AWREADY,
	S0_data0_AXI_WDATA,
	S0_data0_AXI_WSTRB,
	S0_data0_AXI_WVALID,
	S0_data0_AXI_WREADY,
	S0_data0_AXI_BRESP,
	S0_data0_AXI_BVALID,
	S0_data0_AXI_BREADY,
	S0_data0_AXI_ARADDR,
	S0_data0_AXI_ARVALID,
	S0_data0_AXI_ARREADY,
	S0_data0_AXI_RDATA,
	S0_data0_AXI_RRESP,
	S0_data0_AXI_RVALID,
	S0_data0_AXI_RREADY,
	// data1 AXI port
	S0_data1_AXI_ACLK,
	S0_data1_AXI_ARESETN,
	S0_data1_AXI_AWADDR,
	S0_data1_AXI_AWVALID,
	S0_data1_AXI_AWREADY,
	S0_data1_AXI_WDATA,
	S0_data1_AXI_WSTRB,
	S0_data1_AXI_WVALID,
	S0_data1_AXI_WREADY,
	S0_data1_AXI_BRESP,
	S0_data1_AXI_BVALID,
	S0_data1_AXI_BREADY,
	S0_data1_AXI_ARADDR,
	S0_data1_AXI_ARVALID,
	S0_data1_AXI_ARREADY,
	S0_data1_AXI_RDATA,
	S0_data1_AXI_RRESP,
	S0_data1_AXI_RVALID,
	S0_data1_AXI_RREADY,
	// data2 AXI port
	S0_data2_AXI_ACLK,
	S0_data2_AXI_ARESETN,
	S0_data2_AXI_AWADDR,
	S0_data2_AXI_AWVALID,
	S0_data2_AXI_AWREADY,
	S0_data2_AXI_WDATA,
	S0_data2_AXI_WSTRB,
	S0_data2_AXI_WVALID,
	S0_data2_AXI_WREADY,
	S0_data2_AXI_BRESP,
	S0_data2_AXI_BVALID,
	S0_data2_AXI_BREADY,
	S0_data2_AXI_ARADDR,
	S0_data2_AXI_ARVALID,
	S0_data2_AXI_ARREADY,
	S0_data2_AXI_RDATA,
	S0_data2_AXI_RRESP,
	S0_data2_AXI_RVALID,
	S0_data2_AXI_RREADY,
	// data_fixed AXI port
	S1_data_fixed_AXI_ACLK,
	S1_data_fixed_AXI_ARESETN,
	S1_data_fixed_AXI_AWADDR,
	S1_data_fixed_AXI_AWVALID,
	S1_data_fixed_AXI_AWREADY,
	S1_data_fixed_AXI_WDATA,
	S1_data_fixed_AXI_WSTRB,
	S1_data_fixed_AXI_WVALID,
	S1_data_fixed_AXI_WREADY,
	S1_data_fixed_AXI_BRESP,
	S1_data_fixed_AXI_BVALID,
	S1_data_fixed_AXI_BREADY,
	S1_data_fixed_AXI_ARADDR,
	S1_data_fixed_AXI_ARVALID,
	S1_data_fixed_AXI_ARREADY,
	S1_data_fixed_AXI_RDATA,
	S1_data_fixed_AXI_RRESP,
	S1_data_fixed_AXI_RVALID,
	S1_data_fixed_AXI_RREADY,
	// Interrupt lines
	Interrupt_0,
	Interrupt_ctrl0,
	Interrupt_1,
	Interrupt_ctrl1,
	Interrupt_2,
	Interrupt_ctrl2,
	Interrupt_fixed,
	Interrupt_ctrl_fixed,
	busy0,
	busy1,
	busy2,
	busy3,
	busy4,
	busy5,
	busy6,
	busy7,
	//tmp output for verification
	state_reg_out,
	S0_data_AXI_WDATA,
	S0_data_AXI_RDATA,	

);
wire clk;
wire aresetn;
assign clk = S_CLK;
assign aresetn = S_ARESETN;
wire [7:0] owner_id;
assign owner_id = state_reg_out[31:24];

reg reset_latched;
  reg init = 1;
  always @(posedge clk) begin
    if (init) assume (!aresetn);
    if (aresetn) begin    
	case(owner_id)
		`ID0: begin
			assert( S0_data_AXI_WDATA == S0_data0_AXI_WDATA);
			assert( S0_data_AXI_RDATA == S0_data0_AXI_RDATA);
		end
		`ID1: begin
			assert( S0_data_AXI_WDATA == S0_data1_AXI_WDATA);
			assert( S0_data_AXI_RDATA == S0_data1_AXI_RDATA);
		end
		`ID2: begin
			assert( S0_data_AXI_WDATA == S0_data2_AXI_WDATA);
			assert( S0_data_AXI_RDATA == S0_data2_AXI_RDATA);
		end
	endcase
		
    end
    init <= 0;
  end

endmodule
